
module mac ( activ, weight, prev_mac_o, out );
  input [7:0] activ;
  input [7:0] weight;
  input [23:0] prev_mac_o;
  output [23:0] out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003;

  NAND2_X1 U1 ( .A1(n1), .A2(n2), .ZN(out[9]) );
  NAND2_X1 U2 ( .A1(n3), .A2(n4), .ZN(n2) );
  NOR2_X1 U3 ( .A1(n5), .A2(n6), .ZN(n3) );
  NOR2_X1 U4 ( .A1(prev_mac_o[9]), .A2(n7), .ZN(n6) );
  NOR2_X1 U5 ( .A1(n8), .A2(n9), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n10), .A2(n11), .ZN(n1) );
  NAND2_X1 U7 ( .A1(n12), .A2(n13), .ZN(n10) );
  NAND2_X1 U8 ( .A1(prev_mac_o[9]), .A2(n7), .ZN(n13) );
  NAND2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n12) );
  INV_X1 U10 ( .I(prev_mac_o[9]), .ZN(n9) );
  NAND2_X1 U11 ( .A1(n14), .A2(n15), .ZN(out[8]) );
  NAND2_X1 U12 ( .A1(n16), .A2(n17), .ZN(n15) );
  NOR2_X1 U13 ( .A1(n18), .A2(n19), .ZN(n16) );
  NOR2_X1 U14 ( .A1(prev_mac_o[8]), .A2(n20), .ZN(n19) );
  NOR2_X1 U15 ( .A1(n21), .A2(n22), .ZN(n18) );
  NAND2_X1 U16 ( .A1(n23), .A2(n24), .ZN(n14) );
  NAND2_X1 U17 ( .A1(n25), .A2(n26), .ZN(n23) );
  NAND2_X1 U18 ( .A1(n20), .A2(prev_mac_o[8]), .ZN(n26) );
  NAND2_X1 U19 ( .A1(n22), .A2(n21), .ZN(n25) );
  INV_X1 U20 ( .I(prev_mac_o[8]), .ZN(n21) );
  NAND2_X1 U21 ( .A1(n27), .A2(n28), .ZN(out[7]) );
  NAND2_X1 U22 ( .A1(n29), .A2(n30), .ZN(n28) );
  NOR2_X1 U23 ( .A1(n31), .A2(n32), .ZN(n29) );
  NOR2_X1 U24 ( .A1(prev_mac_o[7]), .A2(n33), .ZN(n32) );
  NOR2_X1 U25 ( .A1(n34), .A2(n35), .ZN(n31) );
  NAND2_X1 U26 ( .A1(n36), .A2(n37), .ZN(n27) );
  NAND2_X1 U27 ( .A1(n38), .A2(n39), .ZN(n36) );
  NAND2_X1 U28 ( .A1(n33), .A2(prev_mac_o[7]), .ZN(n39) );
  NAND2_X1 U29 ( .A1(n35), .A2(n34), .ZN(n38) );
  INV_X1 U30 ( .I(prev_mac_o[7]), .ZN(n34) );
  NAND2_X1 U31 ( .A1(n40), .A2(n41), .ZN(out[6]) );
  NAND2_X1 U32 ( .A1(n42), .A2(n43), .ZN(n41) );
  NOR2_X1 U33 ( .A1(n44), .A2(n45), .ZN(n42) );
  NOR2_X1 U34 ( .A1(prev_mac_o[6]), .A2(n46), .ZN(n45) );
  NOR2_X1 U35 ( .A1(n47), .A2(n48), .ZN(n44) );
  NAND2_X1 U36 ( .A1(n49), .A2(n50), .ZN(n40) );
  NAND2_X1 U37 ( .A1(n51), .A2(n52), .ZN(n49) );
  NAND2_X1 U38 ( .A1(n46), .A2(prev_mac_o[6]), .ZN(n52) );
  NAND2_X1 U39 ( .A1(n48), .A2(n47), .ZN(n51) );
  INV_X1 U40 ( .I(prev_mac_o[6]), .ZN(n47) );
  NAND2_X1 U41 ( .A1(n53), .A2(n54), .ZN(out[5]) );
  NAND2_X1 U42 ( .A1(n55), .A2(n56), .ZN(n54) );
  NAND2_X1 U43 ( .A1(n57), .A2(n58), .ZN(n55) );
  NAND2_X1 U44 ( .A1(n59), .A2(prev_mac_o[5]), .ZN(n58) );
  NAND2_X1 U45 ( .A1(n60), .A2(n61), .ZN(n57) );
  NAND2_X1 U46 ( .A1(n62), .A2(n63), .ZN(n53) );
  NOR2_X1 U47 ( .A1(n64), .A2(n65), .ZN(n62) );
  NOR2_X1 U48 ( .A1(prev_mac_o[5]), .A2(n59), .ZN(n65) );
  NOR2_X1 U49 ( .A1(n61), .A2(n60), .ZN(n64) );
  INV_X1 U50 ( .I(prev_mac_o[5]), .ZN(n61) );
  NAND2_X1 U51 ( .A1(n66), .A2(n67), .ZN(out[4]) );
  NAND2_X1 U52 ( .A1(n68), .A2(n69), .ZN(n67) );
  NAND2_X1 U53 ( .A1(n70), .A2(n71), .ZN(n68) );
  NAND2_X1 U54 ( .A1(n72), .A2(prev_mac_o[4]), .ZN(n71) );
  NAND2_X1 U55 ( .A1(n73), .A2(n74), .ZN(n70) );
  NAND2_X1 U56 ( .A1(n75), .A2(n76), .ZN(n66) );
  NOR2_X1 U57 ( .A1(n77), .A2(n78), .ZN(n75) );
  NOR2_X1 U58 ( .A1(prev_mac_o[4]), .A2(n72), .ZN(n78) );
  NOR2_X1 U59 ( .A1(n74), .A2(n73), .ZN(n77) );
  INV_X1 U60 ( .I(prev_mac_o[4]), .ZN(n74) );
  NAND2_X1 U61 ( .A1(n79), .A2(n80), .ZN(out[3]) );
  NAND2_X1 U62 ( .A1(n81), .A2(n82), .ZN(n80) );
  NAND2_X1 U63 ( .A1(n83), .A2(n84), .ZN(n81) );
  NAND2_X1 U64 ( .A1(n85), .A2(prev_mac_o[3]), .ZN(n84) );
  NAND2_X1 U65 ( .A1(n86), .A2(n87), .ZN(n83) );
  NAND2_X1 U66 ( .A1(n88), .A2(n89), .ZN(n79) );
  NOR2_X1 U67 ( .A1(n90), .A2(n91), .ZN(n88) );
  NOR2_X1 U68 ( .A1(prev_mac_o[3]), .A2(n85), .ZN(n91) );
  NOR2_X1 U69 ( .A1(n87), .A2(n86), .ZN(n90) );
  INV_X1 U70 ( .I(prev_mac_o[3]), .ZN(n87) );
  NAND2_X1 U71 ( .A1(n92), .A2(n93), .ZN(out[2]) );
  NAND2_X1 U72 ( .A1(n94), .A2(n95), .ZN(n93) );
  NOR2_X1 U73 ( .A1(n96), .A2(n97), .ZN(n94) );
  NOR2_X1 U74 ( .A1(prev_mac_o[2]), .A2(n98), .ZN(n97) );
  NOR2_X1 U75 ( .A1(n99), .A2(n100), .ZN(n96) );
  NAND2_X1 U76 ( .A1(n101), .A2(n102), .ZN(n92) );
  NAND2_X1 U77 ( .A1(n103), .A2(n104), .ZN(n101) );
  NAND2_X1 U78 ( .A1(n98), .A2(prev_mac_o[2]), .ZN(n104) );
  NAND2_X1 U79 ( .A1(n100), .A2(n99), .ZN(n103) );
  INV_X1 U80 ( .I(prev_mac_o[2]), .ZN(n99) );
  NAND2_X1 U81 ( .A1(n105), .A2(n106), .ZN(out[23]) );
  NAND2_X1 U82 ( .A1(prev_mac_o[23]), .A2(n107), .ZN(n106) );
  INV_X1 U83 ( .I(n108), .ZN(n105) );
  NOR2_X1 U84 ( .A1(n107), .A2(prev_mac_o[23]), .ZN(n108) );
  NAND2_X1 U85 ( .A1(prev_mac_o[22]), .A2(n109), .ZN(n107) );
  INV_X1 U86 ( .I(n110), .ZN(n109) );
  NAND2_X1 U87 ( .A1(n111), .A2(n112), .ZN(out[22]) );
  NAND2_X1 U88 ( .A1(prev_mac_o[22]), .A2(n110), .ZN(n112) );
  INV_X1 U89 ( .I(n113), .ZN(n111) );
  NOR2_X1 U90 ( .A1(n110), .A2(prev_mac_o[22]), .ZN(n113) );
  NAND2_X1 U91 ( .A1(prev_mac_o[21]), .A2(n114), .ZN(n110) );
  NAND2_X1 U92 ( .A1(n115), .A2(n116), .ZN(out[21]) );
  NAND2_X1 U93 ( .A1(prev_mac_o[21]), .A2(n117), .ZN(n116) );
  INV_X1 U94 ( .I(n118), .ZN(n115) );
  NOR2_X1 U95 ( .A1(n117), .A2(prev_mac_o[21]), .ZN(n118) );
  INV_X1 U96 ( .I(n114), .ZN(n117) );
  NOR2_X1 U97 ( .A1(n119), .A2(n120), .ZN(n114) );
  INV_X1 U98 ( .I(prev_mac_o[20]), .ZN(n119) );
  NAND2_X1 U99 ( .A1(n121), .A2(n122), .ZN(out[20]) );
  NAND2_X1 U100 ( .A1(prev_mac_o[20]), .A2(n120), .ZN(n122) );
  INV_X1 U101 ( .I(n123), .ZN(n121) );
  NOR2_X1 U102 ( .A1(n120), .A2(prev_mac_o[20]), .ZN(n123) );
  NAND2_X1 U103 ( .A1(prev_mac_o[19]), .A2(n124), .ZN(n120) );
  NAND2_X1 U104 ( .A1(n125), .A2(n126), .ZN(out[1]) );
  INV_X1 U105 ( .I(n127), .ZN(n126) );
  NOR2_X1 U106 ( .A1(n128), .A2(n129), .ZN(n127) );
  NAND2_X1 U107 ( .A1(n129), .A2(n128), .ZN(n125) );
  NAND2_X1 U108 ( .A1(n130), .A2(n131), .ZN(n129) );
  NAND2_X1 U109 ( .A1(prev_mac_o[1]), .A2(n132), .ZN(n131) );
  INV_X1 U110 ( .I(n133), .ZN(n130) );
  NOR2_X1 U111 ( .A1(n132), .A2(prev_mac_o[1]), .ZN(n133) );
  NAND2_X1 U112 ( .A1(n134), .A2(n135), .ZN(out[19]) );
  NAND2_X1 U113 ( .A1(prev_mac_o[19]), .A2(n136), .ZN(n135) );
  INV_X1 U114 ( .I(n137), .ZN(n134) );
  NOR2_X1 U115 ( .A1(n136), .A2(prev_mac_o[19]), .ZN(n137) );
  INV_X1 U116 ( .I(n124), .ZN(n136) );
  NOR2_X1 U117 ( .A1(n138), .A2(n139), .ZN(n124) );
  INV_X1 U118 ( .I(prev_mac_o[18]), .ZN(n138) );
  NAND2_X1 U119 ( .A1(n140), .A2(n141), .ZN(out[18]) );
  NAND2_X1 U120 ( .A1(prev_mac_o[18]), .A2(n139), .ZN(n141) );
  INV_X1 U121 ( .I(n142), .ZN(n140) );
  NOR2_X1 U122 ( .A1(n139), .A2(prev_mac_o[18]), .ZN(n142) );
  NAND2_X1 U123 ( .A1(prev_mac_o[17]), .A2(n143), .ZN(n139) );
  NAND2_X1 U124 ( .A1(n144), .A2(n145), .ZN(out[17]) );
  NAND2_X1 U125 ( .A1(prev_mac_o[17]), .A2(n146), .ZN(n145) );
  INV_X1 U126 ( .I(n147), .ZN(n144) );
  NOR2_X1 U127 ( .A1(n146), .A2(prev_mac_o[17]), .ZN(n147) );
  NOR2_X1 U128 ( .A1(n143), .A2(n148), .ZN(out[16]) );
  NOR2_X1 U129 ( .A1(prev_mac_o[16]), .A2(n149), .ZN(n148) );
  INV_X1 U130 ( .I(n146), .ZN(n143) );
  NAND2_X1 U131 ( .A1(n149), .A2(prev_mac_o[16]), .ZN(n146) );
  NAND2_X1 U132 ( .A1(n150), .A2(n151), .ZN(n149) );
  NAND2_X1 U133 ( .A1(prev_mac_o[15]), .A2(n152), .ZN(n151) );
  NAND2_X1 U134 ( .A1(n153), .A2(n154), .ZN(n152) );
  NAND2_X1 U135 ( .A1(n155), .A2(n156), .ZN(n150) );
  NAND2_X1 U136 ( .A1(n157), .A2(n158), .ZN(out[15]) );
  NAND2_X1 U137 ( .A1(n159), .A2(n156), .ZN(n158) );
  NAND2_X1 U138 ( .A1(n160), .A2(n161), .ZN(n159) );
  NAND2_X1 U139 ( .A1(prev_mac_o[15]), .A2(n155), .ZN(n161) );
  NAND2_X1 U140 ( .A1(n154), .A2(n162), .ZN(n160) );
  NAND2_X1 U141 ( .A1(n163), .A2(n153), .ZN(n157) );
  INV_X1 U142 ( .I(n156), .ZN(n153) );
  NAND2_X1 U143 ( .A1(n164), .A2(n165), .ZN(n156) );
  NAND2_X1 U144 ( .A1(prev_mac_o[14]), .A2(n166), .ZN(n165) );
  NAND2_X1 U145 ( .A1(n167), .A2(n168), .ZN(n166) );
  NAND2_X1 U146 ( .A1(n169), .A2(n170), .ZN(n164) );
  NOR2_X1 U147 ( .A1(n171), .A2(n172), .ZN(n163) );
  NOR2_X1 U148 ( .A1(prev_mac_o[15]), .A2(n155), .ZN(n172) );
  NOR2_X1 U149 ( .A1(n154), .A2(n162), .ZN(n171) );
  INV_X1 U150 ( .I(prev_mac_o[15]), .ZN(n162) );
  INV_X1 U151 ( .I(n155), .ZN(n154) );
  NAND2_X1 U152 ( .A1(n173), .A2(n174), .ZN(n155) );
  NAND2_X1 U153 ( .A1(n175), .A2(n176), .ZN(n174) );
  NOR2_X1 U154 ( .A1(n177), .A2(n178), .ZN(n173) );
  INV_X1 U155 ( .I(n179), .ZN(n177) );
  NAND2_X1 U156 ( .A1(n180), .A2(n181), .ZN(out[14]) );
  NAND2_X1 U157 ( .A1(n182), .A2(n170), .ZN(n181) );
  NAND2_X1 U158 ( .A1(n183), .A2(n184), .ZN(n182) );
  NAND2_X1 U159 ( .A1(n169), .A2(prev_mac_o[14]), .ZN(n184) );
  NAND2_X1 U160 ( .A1(n168), .A2(n185), .ZN(n183) );
  NAND2_X1 U161 ( .A1(n186), .A2(n167), .ZN(n180) );
  INV_X1 U162 ( .I(n170), .ZN(n167) );
  NAND2_X1 U163 ( .A1(n187), .A2(n188), .ZN(n170) );
  NAND2_X1 U164 ( .A1(prev_mac_o[13]), .A2(n189), .ZN(n188) );
  NAND2_X1 U165 ( .A1(n190), .A2(n191), .ZN(n189) );
  NAND2_X1 U166 ( .A1(n192), .A2(n193), .ZN(n187) );
  NOR2_X1 U167 ( .A1(n194), .A2(n195), .ZN(n186) );
  NOR2_X1 U168 ( .A1(prev_mac_o[14]), .A2(n169), .ZN(n195) );
  INV_X1 U169 ( .I(n168), .ZN(n169) );
  NOR2_X1 U170 ( .A1(n185), .A2(n168), .ZN(n194) );
  NAND2_X1 U171 ( .A1(n196), .A2(n197), .ZN(n168) );
  NAND2_X1 U172 ( .A1(n198), .A2(n175), .ZN(n197) );
  INV_X1 U173 ( .I(n199), .ZN(n196) );
  NOR2_X1 U174 ( .A1(n175), .A2(n198), .ZN(n199) );
  NOR2_X1 U175 ( .A1(n200), .A2(n178), .ZN(n198) );
  NOR2_X1 U176 ( .A1(n201), .A2(n202), .ZN(n178) );
  INV_X1 U177 ( .I(n176), .ZN(n200) );
  NAND2_X1 U178 ( .A1(n202), .A2(n201), .ZN(n176) );
  NAND2_X1 U179 ( .A1(n203), .A2(n204), .ZN(n201) );
  NAND2_X1 U180 ( .A1(n205), .A2(n179), .ZN(n202) );
  NAND2_X1 U181 ( .A1(activ[7]), .A2(n206), .ZN(n179) );
  NAND2_X1 U182 ( .A1(n207), .A2(n208), .ZN(n205) );
  NAND2_X1 U183 ( .A1(activ[7]), .A2(weight[7]), .ZN(n208) );
  INV_X1 U184 ( .I(n206), .ZN(n207) );
  NAND2_X1 U185 ( .A1(n209), .A2(n210), .ZN(n206) );
  NAND2_X1 U186 ( .A1(n211), .A2(n212), .ZN(n210) );
  NAND2_X1 U187 ( .A1(n213), .A2(n214), .ZN(n211) );
  NAND2_X1 U188 ( .A1(n215), .A2(n216), .ZN(n209) );
  NAND2_X1 U189 ( .A1(n217), .A2(n218), .ZN(n175) );
  NAND2_X1 U190 ( .A1(n219), .A2(n220), .ZN(n218) );
  INV_X1 U191 ( .I(prev_mac_o[14]), .ZN(n185) );
  NAND2_X1 U192 ( .A1(n221), .A2(n222), .ZN(out[13]) );
  NAND2_X1 U193 ( .A1(n223), .A2(n193), .ZN(n222) );
  NAND2_X1 U194 ( .A1(n224), .A2(n225), .ZN(n223) );
  NAND2_X1 U195 ( .A1(n192), .A2(prev_mac_o[13]), .ZN(n225) );
  NAND2_X1 U196 ( .A1(n191), .A2(n226), .ZN(n224) );
  NAND2_X1 U197 ( .A1(n227), .A2(n190), .ZN(n221) );
  INV_X1 U198 ( .I(n193), .ZN(n190) );
  NAND2_X1 U199 ( .A1(n228), .A2(n229), .ZN(n193) );
  NAND2_X1 U200 ( .A1(prev_mac_o[12]), .A2(n230), .ZN(n229) );
  NAND2_X1 U201 ( .A1(n231), .A2(n232), .ZN(n230) );
  NAND2_X1 U202 ( .A1(n233), .A2(n234), .ZN(n228) );
  NOR2_X1 U203 ( .A1(n235), .A2(n236), .ZN(n227) );
  NOR2_X1 U204 ( .A1(prev_mac_o[13]), .A2(n192), .ZN(n236) );
  INV_X1 U205 ( .I(n191), .ZN(n192) );
  NOR2_X1 U206 ( .A1(n226), .A2(n191), .ZN(n235) );
  NAND2_X1 U207 ( .A1(n237), .A2(n238), .ZN(n191) );
  NAND2_X1 U208 ( .A1(n239), .A2(n219), .ZN(n238) );
  INV_X1 U209 ( .I(n240), .ZN(n239) );
  NAND2_X1 U210 ( .A1(n241), .A2(n240), .ZN(n237) );
  NAND2_X1 U211 ( .A1(n220), .A2(n217), .ZN(n240) );
  NAND2_X1 U212 ( .A1(n242), .A2(n243), .ZN(n217) );
  NAND2_X1 U213 ( .A1(n244), .A2(n245), .ZN(n243) );
  NAND2_X1 U214 ( .A1(n246), .A2(n203), .ZN(n245) );
  NAND2_X1 U215 ( .A1(n247), .A2(n204), .ZN(n244) );
  NAND2_X1 U216 ( .A1(n248), .A2(n249), .ZN(n220) );
  NOR2_X1 U217 ( .A1(n250), .A2(n251), .ZN(n248) );
  NOR2_X1 U218 ( .A1(n246), .A2(n203), .ZN(n251) );
  INV_X1 U219 ( .I(n247), .ZN(n203) );
  INV_X1 U220 ( .I(n204), .ZN(n246) );
  NOR2_X1 U221 ( .A1(n247), .A2(n204), .ZN(n250) );
  NAND2_X1 U222 ( .A1(n252), .A2(n253), .ZN(n204) );
  NAND2_X1 U223 ( .A1(n254), .A2(n255), .ZN(n253) );
  NAND2_X1 U224 ( .A1(n256), .A2(n257), .ZN(n254) );
  NAND2_X1 U225 ( .A1(n258), .A2(n259), .ZN(n252) );
  NAND2_X1 U226 ( .A1(n260), .A2(n261), .ZN(n247) );
  INV_X1 U227 ( .I(n262), .ZN(n261) );
  NOR2_X1 U228 ( .A1(n212), .A2(n263), .ZN(n262) );
  NAND2_X1 U229 ( .A1(n263), .A2(n212), .ZN(n260) );
  NAND2_X1 U230 ( .A1(n264), .A2(n265), .ZN(n212) );
  NAND2_X1 U231 ( .A1(n266), .A2(n267), .ZN(n265) );
  NAND2_X1 U232 ( .A1(n268), .A2(n269), .ZN(n266) );
  NAND2_X1 U233 ( .A1(n270), .A2(n271), .ZN(n264) );
  NAND2_X1 U234 ( .A1(n272), .A2(n273), .ZN(n263) );
  NAND2_X1 U235 ( .A1(n216), .A2(n214), .ZN(n273) );
  INV_X1 U236 ( .I(n213), .ZN(n216) );
  NAND2_X1 U237 ( .A1(n215), .A2(n213), .ZN(n272) );
  NAND2_X1 U238 ( .A1(activ[7]), .A2(weight[6]), .ZN(n213) );
  INV_X1 U239 ( .I(n214), .ZN(n215) );
  NAND2_X1 U240 ( .A1(weight[7]), .A2(activ[6]), .ZN(n214) );
  INV_X1 U241 ( .I(n219), .ZN(n241) );
  NAND2_X1 U242 ( .A1(n274), .A2(n275), .ZN(n219) );
  INV_X1 U243 ( .I(prev_mac_o[13]), .ZN(n226) );
  NAND2_X1 U244 ( .A1(n276), .A2(n277), .ZN(out[12]) );
  NAND2_X1 U245 ( .A1(n278), .A2(n234), .ZN(n277) );
  NAND2_X1 U246 ( .A1(n279), .A2(n280), .ZN(n278) );
  NAND2_X1 U247 ( .A1(n233), .A2(prev_mac_o[12]), .ZN(n280) );
  NAND2_X1 U248 ( .A1(n232), .A2(n281), .ZN(n279) );
  NAND2_X1 U249 ( .A1(n282), .A2(n231), .ZN(n276) );
  INV_X1 U250 ( .I(n234), .ZN(n231) );
  NAND2_X1 U251 ( .A1(n283), .A2(n284), .ZN(n234) );
  NAND2_X1 U252 ( .A1(prev_mac_o[11]), .A2(n285), .ZN(n284) );
  NAND2_X1 U253 ( .A1(n286), .A2(n287), .ZN(n285) );
  NAND2_X1 U254 ( .A1(n288), .A2(n289), .ZN(n283) );
  NOR2_X1 U255 ( .A1(n290), .A2(n291), .ZN(n282) );
  NOR2_X1 U256 ( .A1(prev_mac_o[12]), .A2(n233), .ZN(n291) );
  INV_X1 U257 ( .I(n232), .ZN(n233) );
  NOR2_X1 U258 ( .A1(n281), .A2(n232), .ZN(n290) );
  NAND2_X1 U259 ( .A1(n275), .A2(n292), .ZN(n232) );
  NAND2_X1 U260 ( .A1(n293), .A2(n294), .ZN(n292) );
  NAND2_X1 U261 ( .A1(n295), .A2(n274), .ZN(n294) );
  NAND2_X1 U262 ( .A1(n296), .A2(n297), .ZN(n274) );
  INV_X1 U263 ( .I(n298), .ZN(n293) );
  NAND2_X1 U264 ( .A1(n295), .A2(n298), .ZN(n275) );
  NAND2_X1 U265 ( .A1(n299), .A2(n300), .ZN(n298) );
  NAND2_X1 U266 ( .A1(n301), .A2(n302), .ZN(n300) );
  INV_X1 U267 ( .I(n303), .ZN(n295) );
  NOR2_X1 U268 ( .A1(n296), .A2(n297), .ZN(n303) );
  INV_X1 U269 ( .I(n304), .ZN(n297) );
  NAND2_X1 U270 ( .A1(n249), .A2(n305), .ZN(n304) );
  NAND2_X1 U271 ( .A1(n306), .A2(n307), .ZN(n305) );
  INV_X1 U272 ( .I(n242), .ZN(n249) );
  NOR2_X1 U273 ( .A1(n307), .A2(n306), .ZN(n242) );
  NOR2_X1 U274 ( .A1(n308), .A2(n309), .ZN(n306) );
  INV_X1 U275 ( .I(n310), .ZN(n309) );
  NAND2_X1 U276 ( .A1(n256), .A2(n311), .ZN(n310) );
  NOR2_X1 U277 ( .A1(n311), .A2(n256), .ZN(n308) );
  INV_X1 U278 ( .I(n258), .ZN(n256) );
  NOR2_X1 U279 ( .A1(n312), .A2(n313), .ZN(n258) );
  NOR2_X1 U280 ( .A1(n267), .A2(n314), .ZN(n313) );
  INV_X1 U281 ( .I(n315), .ZN(n312) );
  NAND2_X1 U282 ( .A1(n314), .A2(n267), .ZN(n315) );
  NAND2_X1 U283 ( .A1(n316), .A2(n317), .ZN(n267) );
  NAND2_X1 U284 ( .A1(n318), .A2(n319), .ZN(n317) );
  NAND2_X1 U285 ( .A1(n320), .A2(n321), .ZN(n318) );
  NAND2_X1 U286 ( .A1(n322), .A2(n323), .ZN(n316) );
  NAND2_X1 U287 ( .A1(n324), .A2(n325), .ZN(n314) );
  NAND2_X1 U288 ( .A1(n271), .A2(n269), .ZN(n325) );
  INV_X1 U289 ( .I(n268), .ZN(n271) );
  NAND2_X1 U290 ( .A1(n270), .A2(n268), .ZN(n324) );
  NAND2_X1 U291 ( .A1(weight[6]), .A2(activ[6]), .ZN(n268) );
  INV_X1 U292 ( .I(n269), .ZN(n270) );
  NAND2_X1 U293 ( .A1(weight[7]), .A2(activ[5]), .ZN(n269) );
  NOR2_X1 U294 ( .A1(n326), .A2(n327), .ZN(n311) );
  INV_X1 U295 ( .I(n328), .ZN(n327) );
  NAND2_X1 U296 ( .A1(n259), .A2(n255), .ZN(n328) );
  NOR2_X1 U297 ( .A1(n255), .A2(n259), .ZN(n326) );
  INV_X1 U298 ( .I(n257), .ZN(n259) );
  NAND2_X1 U299 ( .A1(activ[7]), .A2(weight[5]), .ZN(n257) );
  NAND2_X1 U300 ( .A1(n329), .A2(n330), .ZN(n255) );
  NAND2_X1 U301 ( .A1(n331), .A2(n332), .ZN(n330) );
  NAND2_X1 U302 ( .A1(n333), .A2(n334), .ZN(n307) );
  NAND2_X1 U303 ( .A1(n335), .A2(n336), .ZN(n334) );
  NAND2_X1 U304 ( .A1(n337), .A2(n338), .ZN(n335) );
  INV_X1 U305 ( .I(n339), .ZN(n333) );
  NOR2_X1 U306 ( .A1(n337), .A2(n338), .ZN(n339) );
  INV_X1 U307 ( .I(prev_mac_o[12]), .ZN(n281) );
  NAND2_X1 U308 ( .A1(n340), .A2(n341), .ZN(out[11]) );
  NAND2_X1 U309 ( .A1(n342), .A2(n289), .ZN(n341) );
  NAND2_X1 U310 ( .A1(n343), .A2(n344), .ZN(n342) );
  NAND2_X1 U311 ( .A1(n288), .A2(prev_mac_o[11]), .ZN(n344) );
  NAND2_X1 U312 ( .A1(n287), .A2(n345), .ZN(n343) );
  NAND2_X1 U313 ( .A1(n346), .A2(n286), .ZN(n340) );
  INV_X1 U314 ( .I(n289), .ZN(n286) );
  NAND2_X1 U315 ( .A1(n347), .A2(n348), .ZN(n289) );
  NAND2_X1 U316 ( .A1(prev_mac_o[10]), .A2(n349), .ZN(n348) );
  NAND2_X1 U317 ( .A1(n350), .A2(n351), .ZN(n349) );
  NAND2_X1 U318 ( .A1(n352), .A2(n353), .ZN(n347) );
  NOR2_X1 U319 ( .A1(n354), .A2(n355), .ZN(n346) );
  NOR2_X1 U320 ( .A1(prev_mac_o[11]), .A2(n288), .ZN(n355) );
  INV_X1 U321 ( .I(n287), .ZN(n288) );
  NOR2_X1 U322 ( .A1(n345), .A2(n287), .ZN(n354) );
  NAND2_X1 U323 ( .A1(n356), .A2(n357), .ZN(n287) );
  NAND2_X1 U324 ( .A1(n358), .A2(n301), .ZN(n357) );
  INV_X1 U325 ( .I(n359), .ZN(n358) );
  NAND2_X1 U326 ( .A1(n360), .A2(n359), .ZN(n356) );
  NAND2_X1 U327 ( .A1(n302), .A2(n299), .ZN(n359) );
  NAND2_X1 U328 ( .A1(n361), .A2(n362), .ZN(n299) );
  NOR2_X1 U329 ( .A1(n296), .A2(n363), .ZN(n361) );
  NOR2_X1 U330 ( .A1(n364), .A2(n365), .ZN(n363) );
  NOR2_X1 U331 ( .A1(n366), .A2(n367), .ZN(n296) );
  NAND2_X1 U332 ( .A1(n368), .A2(n369), .ZN(n302) );
  NOR2_X1 U333 ( .A1(n370), .A2(n371), .ZN(n368) );
  NOR2_X1 U334 ( .A1(n367), .A2(n364), .ZN(n371) );
  INV_X1 U335 ( .I(n366), .ZN(n364) );
  INV_X1 U336 ( .I(n365), .ZN(n367) );
  NOR2_X1 U337 ( .A1(n365), .A2(n366), .ZN(n370) );
  NAND2_X1 U338 ( .A1(n372), .A2(n373), .ZN(n366) );
  INV_X1 U339 ( .I(n374), .ZN(n373) );
  NOR2_X1 U340 ( .A1(n337), .A2(n375), .ZN(n374) );
  NAND2_X1 U341 ( .A1(n375), .A2(n337), .ZN(n372) );
  NOR2_X1 U342 ( .A1(n376), .A2(n377), .ZN(n337) );
  NOR2_X1 U343 ( .A1(n378), .A2(n379), .ZN(n377) );
  NOR2_X1 U344 ( .A1(n331), .A2(n380), .ZN(n376) );
  INV_X1 U345 ( .I(n378), .ZN(n380) );
  NAND2_X1 U346 ( .A1(n329), .A2(n332), .ZN(n378) );
  NAND2_X1 U347 ( .A1(n381), .A2(n382), .ZN(n332) );
  NAND2_X1 U348 ( .A1(activ[6]), .A2(weight[5]), .ZN(n382) );
  INV_X1 U349 ( .I(n383), .ZN(n381) );
  NAND2_X1 U350 ( .A1(activ[6]), .A2(n383), .ZN(n329) );
  NAND2_X1 U351 ( .A1(n384), .A2(n385), .ZN(n383) );
  NAND2_X1 U352 ( .A1(n386), .A2(n387), .ZN(n385) );
  NOR2_X1 U353 ( .A1(n388), .A2(n389), .ZN(n386) );
  NOR2_X1 U354 ( .A1(n390), .A2(n391), .ZN(n384) );
  NOR2_X1 U355 ( .A1(n392), .A2(n393), .ZN(n391) );
  INV_X1 U356 ( .I(n379), .ZN(n331) );
  NAND2_X1 U357 ( .A1(n394), .A2(n395), .ZN(n379) );
  INV_X1 U358 ( .I(n396), .ZN(n395) );
  NOR2_X1 U359 ( .A1(n319), .A2(n397), .ZN(n396) );
  NAND2_X1 U360 ( .A1(n397), .A2(n319), .ZN(n394) );
  NAND2_X1 U361 ( .A1(n398), .A2(n399), .ZN(n319) );
  NAND2_X1 U362 ( .A1(n400), .A2(n401), .ZN(n399) );
  NAND2_X1 U363 ( .A1(n402), .A2(n403), .ZN(n400) );
  NAND2_X1 U364 ( .A1(n404), .A2(n405), .ZN(n398) );
  NAND2_X1 U365 ( .A1(n406), .A2(n407), .ZN(n397) );
  NAND2_X1 U366 ( .A1(n323), .A2(n321), .ZN(n407) );
  NAND2_X1 U367 ( .A1(n322), .A2(n320), .ZN(n406) );
  INV_X1 U368 ( .I(n323), .ZN(n320) );
  NOR2_X1 U369 ( .A1(n408), .A2(n388), .ZN(n323) );
  INV_X1 U370 ( .I(n321), .ZN(n322) );
  NAND2_X1 U371 ( .A1(weight[7]), .A2(activ[4]), .ZN(n321) );
  NAND2_X1 U372 ( .A1(n409), .A2(n410), .ZN(n375) );
  NAND2_X1 U373 ( .A1(n411), .A2(n412), .ZN(n410) );
  NAND2_X1 U374 ( .A1(n338), .A2(n336), .ZN(n409) );
  INV_X1 U375 ( .I(n411), .ZN(n336) );
  NOR2_X1 U376 ( .A1(n413), .A2(n414), .ZN(n411) );
  NOR2_X1 U377 ( .A1(n415), .A2(n416), .ZN(n414) );
  NOR2_X1 U378 ( .A1(n417), .A2(n418), .ZN(n415) );
  INV_X1 U379 ( .I(n419), .ZN(n413) );
  NAND2_X1 U380 ( .A1(n417), .A2(n418), .ZN(n419) );
  INV_X1 U381 ( .I(n412), .ZN(n338) );
  NAND2_X1 U382 ( .A1(activ[7]), .A2(weight[4]), .ZN(n412) );
  NAND2_X1 U383 ( .A1(n420), .A2(n421), .ZN(n365) );
  NAND2_X1 U384 ( .A1(n422), .A2(n423), .ZN(n421) );
  INV_X1 U385 ( .I(n301), .ZN(n360) );
  NAND2_X1 U386 ( .A1(n424), .A2(n425), .ZN(n301) );
  NAND2_X1 U387 ( .A1(n426), .A2(n427), .ZN(n425) );
  INV_X1 U388 ( .I(n428), .ZN(n426) );
  NAND2_X1 U389 ( .A1(n429), .A2(n427), .ZN(n424) );
  INV_X1 U390 ( .I(prev_mac_o[11]), .ZN(n345) );
  NAND2_X1 U391 ( .A1(n430), .A2(n431), .ZN(out[10]) );
  NAND2_X1 U392 ( .A1(n432), .A2(n353), .ZN(n431) );
  NOR2_X1 U393 ( .A1(n433), .A2(n434), .ZN(n432) );
  NOR2_X1 U394 ( .A1(prev_mac_o[10]), .A2(n351), .ZN(n434) );
  NOR2_X1 U395 ( .A1(n435), .A2(n352), .ZN(n433) );
  NAND2_X1 U396 ( .A1(n436), .A2(n350), .ZN(n430) );
  INV_X1 U397 ( .I(n353), .ZN(n350) );
  NAND2_X1 U398 ( .A1(n437), .A2(n438), .ZN(n353) );
  NAND2_X1 U399 ( .A1(prev_mac_o[9]), .A2(n439), .ZN(n438) );
  NAND2_X1 U400 ( .A1(n11), .A2(n7), .ZN(n439) );
  INV_X1 U401 ( .I(n4), .ZN(n11) );
  NAND2_X1 U402 ( .A1(n8), .A2(n4), .ZN(n437) );
  NAND2_X1 U403 ( .A1(n440), .A2(n441), .ZN(n4) );
  NAND2_X1 U404 ( .A1(prev_mac_o[8]), .A2(n442), .ZN(n441) );
  NAND2_X1 U405 ( .A1(n24), .A2(n20), .ZN(n442) );
  INV_X1 U406 ( .I(n22), .ZN(n20) );
  INV_X1 U407 ( .I(n17), .ZN(n24) );
  NAND2_X1 U408 ( .A1(n22), .A2(n17), .ZN(n440) );
  NAND2_X1 U409 ( .A1(n443), .A2(n444), .ZN(n17) );
  NAND2_X1 U410 ( .A1(prev_mac_o[7]), .A2(n445), .ZN(n444) );
  NAND2_X1 U411 ( .A1(n37), .A2(n33), .ZN(n445) );
  INV_X1 U412 ( .I(n30), .ZN(n37) );
  NAND2_X1 U413 ( .A1(n35), .A2(n30), .ZN(n443) );
  NAND2_X1 U414 ( .A1(n446), .A2(n447), .ZN(n30) );
  NAND2_X1 U415 ( .A1(prev_mac_o[6]), .A2(n448), .ZN(n447) );
  NAND2_X1 U416 ( .A1(n50), .A2(n46), .ZN(n448) );
  INV_X1 U417 ( .I(n48), .ZN(n46) );
  INV_X1 U418 ( .I(n43), .ZN(n50) );
  NAND2_X1 U419 ( .A1(n48), .A2(n43), .ZN(n446) );
  NAND2_X1 U420 ( .A1(n449), .A2(n450), .ZN(n43) );
  NAND2_X1 U421 ( .A1(prev_mac_o[5]), .A2(n451), .ZN(n450) );
  NAND2_X1 U422 ( .A1(n63), .A2(n60), .ZN(n451) );
  INV_X1 U423 ( .I(n56), .ZN(n63) );
  NAND2_X1 U424 ( .A1(n59), .A2(n56), .ZN(n449) );
  NAND2_X1 U425 ( .A1(n452), .A2(n453), .ZN(n56) );
  NAND2_X1 U426 ( .A1(prev_mac_o[4]), .A2(n454), .ZN(n453) );
  NAND2_X1 U427 ( .A1(n76), .A2(n73), .ZN(n454) );
  INV_X1 U428 ( .I(n72), .ZN(n73) );
  INV_X1 U429 ( .I(n69), .ZN(n76) );
  NAND2_X1 U430 ( .A1(n72), .A2(n69), .ZN(n452) );
  NAND2_X1 U431 ( .A1(n455), .A2(n456), .ZN(n69) );
  NAND2_X1 U432 ( .A1(prev_mac_o[3]), .A2(n457), .ZN(n456) );
  NAND2_X1 U433 ( .A1(n89), .A2(n86), .ZN(n457) );
  INV_X1 U434 ( .I(n82), .ZN(n89) );
  NAND2_X1 U435 ( .A1(n85), .A2(n82), .ZN(n455) );
  NAND2_X1 U436 ( .A1(n458), .A2(n459), .ZN(n82) );
  NAND2_X1 U437 ( .A1(prev_mac_o[2]), .A2(n460), .ZN(n459) );
  NAND2_X1 U438 ( .A1(n102), .A2(n98), .ZN(n460) );
  INV_X1 U439 ( .I(n100), .ZN(n98) );
  NAND2_X1 U440 ( .A1(n100), .A2(n95), .ZN(n458) );
  INV_X1 U441 ( .I(n102), .ZN(n95) );
  NOR2_X1 U442 ( .A1(n461), .A2(n462), .ZN(n102) );
  INV_X1 U443 ( .I(n463), .ZN(n462) );
  NAND2_X1 U444 ( .A1(prev_mac_o[1]), .A2(n464), .ZN(n463) );
  NAND2_X1 U445 ( .A1(n128), .A2(n132), .ZN(n464) );
  NOR2_X1 U446 ( .A1(n132), .A2(n128), .ZN(n461) );
  NOR2_X1 U447 ( .A1(n465), .A2(n466), .ZN(n128) );
  INV_X1 U448 ( .I(n467), .ZN(n466) );
  NAND2_X1 U449 ( .A1(n468), .A2(n469), .ZN(n467) );
  NOR2_X1 U450 ( .A1(n469), .A2(n468), .ZN(n465) );
  NOR2_X1 U451 ( .A1(n470), .A2(n471), .ZN(n468) );
  NAND2_X1 U452 ( .A1(prev_mac_o[0]), .A2(n472), .ZN(n132) );
  NAND2_X1 U453 ( .A1(n473), .A2(n474), .ZN(n100) );
  NAND2_X1 U454 ( .A1(n475), .A2(n476), .ZN(n474) );
  INV_X1 U455 ( .I(n477), .ZN(n473) );
  NOR2_X1 U456 ( .A1(n476), .A2(n475), .ZN(n477) );
  NOR2_X1 U457 ( .A1(n478), .A2(n479), .ZN(n476) );
  INV_X1 U458 ( .I(n480), .ZN(n479) );
  NAND2_X1 U459 ( .A1(n481), .A2(n482), .ZN(n480) );
  NOR2_X1 U460 ( .A1(n482), .A2(n481), .ZN(n478) );
  NAND2_X1 U461 ( .A1(activ[2]), .A2(weight[0]), .ZN(n482) );
  INV_X1 U462 ( .I(n86), .ZN(n85) );
  NAND2_X1 U463 ( .A1(n483), .A2(n484), .ZN(n86) );
  NAND2_X1 U464 ( .A1(n485), .A2(n486), .ZN(n484) );
  INV_X1 U465 ( .I(n487), .ZN(n486) );
  NAND2_X1 U466 ( .A1(n487), .A2(n488), .ZN(n483) );
  NAND2_X1 U467 ( .A1(n489), .A2(n490), .ZN(n487) );
  NAND2_X1 U468 ( .A1(n491), .A2(n492), .ZN(n490) );
  NAND2_X1 U469 ( .A1(n493), .A2(n494), .ZN(n489) );
  NOR2_X1 U470 ( .A1(n495), .A2(n496), .ZN(n72) );
  INV_X1 U471 ( .I(n497), .ZN(n496) );
  NAND2_X1 U472 ( .A1(n498), .A2(n499), .ZN(n497) );
  NOR2_X1 U473 ( .A1(n499), .A2(n498), .ZN(n495) );
  NOR2_X1 U474 ( .A1(n500), .A2(n501), .ZN(n498) );
  INV_X1 U475 ( .I(n502), .ZN(n501) );
  INV_X1 U476 ( .I(n60), .ZN(n59) );
  NAND2_X1 U477 ( .A1(n503), .A2(n504), .ZN(n60) );
  NAND2_X1 U478 ( .A1(n505), .A2(n506), .ZN(n504) );
  INV_X1 U479 ( .I(n507), .ZN(n505) );
  NAND2_X1 U480 ( .A1(n508), .A2(n507), .ZN(n503) );
  NAND2_X1 U481 ( .A1(n509), .A2(n510), .ZN(n507) );
  NAND2_X1 U482 ( .A1(n511), .A2(n512), .ZN(n48) );
  INV_X1 U483 ( .I(n513), .ZN(n512) );
  NOR2_X1 U484 ( .A1(n514), .A2(n515), .ZN(n513) );
  NAND2_X1 U485 ( .A1(n515), .A2(n514), .ZN(n511) );
  NAND2_X1 U486 ( .A1(n516), .A2(n517), .ZN(n514) );
  INV_X1 U487 ( .I(n33), .ZN(n35) );
  NOR2_X1 U488 ( .A1(n518), .A2(n519), .ZN(n33) );
  NOR2_X1 U489 ( .A1(n520), .A2(n521), .ZN(n519) );
  NOR2_X1 U490 ( .A1(n522), .A2(n523), .ZN(n518) );
  INV_X1 U491 ( .I(n521), .ZN(n522) );
  NAND2_X1 U492 ( .A1(n524), .A2(n525), .ZN(n521) );
  NAND2_X1 U493 ( .A1(n526), .A2(n527), .ZN(n525) );
  NAND2_X1 U494 ( .A1(n528), .A2(n529), .ZN(n524) );
  NAND2_X1 U495 ( .A1(n530), .A2(n531), .ZN(n22) );
  NAND2_X1 U496 ( .A1(n532), .A2(n533), .ZN(n531) );
  NAND2_X1 U497 ( .A1(n534), .A2(n535), .ZN(n530) );
  INV_X1 U498 ( .I(n7), .ZN(n8) );
  NAND2_X1 U499 ( .A1(n536), .A2(n428), .ZN(n7) );
  NAND2_X1 U500 ( .A1(n537), .A2(n538), .ZN(n536) );
  NAND2_X1 U501 ( .A1(n533), .A2(n535), .ZN(n538) );
  INV_X1 U502 ( .I(n532), .ZN(n535) );
  NAND2_X1 U503 ( .A1(n539), .A2(n540), .ZN(n537) );
  NAND2_X1 U504 ( .A1(n541), .A2(n542), .ZN(n540) );
  NAND2_X1 U505 ( .A1(n543), .A2(n544), .ZN(n539) );
  NAND2_X1 U506 ( .A1(n545), .A2(n546), .ZN(n436) );
  NAND2_X1 U507 ( .A1(n351), .A2(prev_mac_o[10]), .ZN(n546) );
  NAND2_X1 U508 ( .A1(n352), .A2(n435), .ZN(n545) );
  INV_X1 U509 ( .I(prev_mac_o[10]), .ZN(n435) );
  INV_X1 U510 ( .I(n351), .ZN(n352) );
  NOR2_X1 U511 ( .A1(n547), .A2(n548), .ZN(n351) );
  NOR2_X1 U512 ( .A1(n549), .A2(n428), .ZN(n548) );
  INV_X1 U513 ( .I(n550), .ZN(n547) );
  NAND2_X1 U514 ( .A1(n549), .A2(n428), .ZN(n550) );
  NAND2_X1 U515 ( .A1(n551), .A2(n552), .ZN(n428) );
  NOR2_X1 U516 ( .A1(n429), .A2(n532), .ZN(n552) );
  NOR2_X1 U517 ( .A1(n553), .A2(n554), .ZN(n532) );
  NOR2_X1 U518 ( .A1(n555), .A2(n528), .ZN(n554) );
  INV_X1 U519 ( .I(n527), .ZN(n528) );
  NAND2_X1 U520 ( .A1(n516), .A2(n556), .ZN(n527) );
  NAND2_X1 U521 ( .A1(n515), .A2(n517), .ZN(n556) );
  NAND2_X1 U522 ( .A1(n557), .A2(n558), .ZN(n517) );
  NAND2_X1 U523 ( .A1(activ[6]), .A2(weight[0]), .ZN(n558) );
  INV_X1 U524 ( .I(n559), .ZN(n557) );
  NAND2_X1 U525 ( .A1(n560), .A2(n561), .ZN(n515) );
  NAND2_X1 U526 ( .A1(n562), .A2(n563), .ZN(n561) );
  INV_X1 U527 ( .I(n564), .ZN(n560) );
  NOR2_X1 U528 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U529 ( .A1(n565), .A2(n566), .ZN(n562) );
  NOR2_X1 U530 ( .A1(n567), .A2(n568), .ZN(n565) );
  NOR2_X1 U531 ( .A1(n388), .A2(n569), .ZN(n568) );
  NAND2_X1 U532 ( .A1(activ[6]), .A2(n559), .ZN(n516) );
  NAND2_X1 U533 ( .A1(n510), .A2(n570), .ZN(n559) );
  NAND2_X1 U534 ( .A1(n506), .A2(n509), .ZN(n570) );
  NAND2_X1 U535 ( .A1(n571), .A2(n572), .ZN(n509) );
  NAND2_X1 U536 ( .A1(activ[5]), .A2(weight[0]), .ZN(n572) );
  INV_X1 U537 ( .I(n508), .ZN(n506) );
  NAND2_X1 U538 ( .A1(n573), .A2(n574), .ZN(n508) );
  INV_X1 U539 ( .I(n575), .ZN(n574) );
  NOR2_X1 U540 ( .A1(n576), .A2(n577), .ZN(n575) );
  NAND2_X1 U541 ( .A1(n577), .A2(n576), .ZN(n573) );
  NAND2_X1 U542 ( .A1(n578), .A2(n579), .ZN(n577) );
  NAND2_X1 U543 ( .A1(n580), .A2(n581), .ZN(n579) );
  INV_X1 U544 ( .I(n582), .ZN(n578) );
  NOR2_X1 U545 ( .A1(n581), .A2(n580), .ZN(n582) );
  INV_X1 U546 ( .I(n583), .ZN(n580) );
  NAND2_X1 U547 ( .A1(activ[5]), .A2(n584), .ZN(n510) );
  INV_X1 U548 ( .I(n571), .ZN(n584) );
  NOR2_X1 U549 ( .A1(n500), .A2(n585), .ZN(n571) );
  INV_X1 U550 ( .I(n586), .ZN(n585) );
  NAND2_X1 U551 ( .A1(n499), .A2(n502), .ZN(n586) );
  NAND2_X1 U552 ( .A1(n587), .A2(n588), .ZN(n502) );
  NOR2_X1 U553 ( .A1(n589), .A2(n590), .ZN(n499) );
  INV_X1 U554 ( .I(n591), .ZN(n590) );
  NAND2_X1 U555 ( .A1(n592), .A2(n593), .ZN(n591) );
  NOR2_X1 U556 ( .A1(n593), .A2(n592), .ZN(n589) );
  NOR2_X1 U557 ( .A1(n594), .A2(n595), .ZN(n593) );
  NOR2_X1 U558 ( .A1(n596), .A2(n597), .ZN(n595) );
  NOR2_X1 U559 ( .A1(n598), .A2(n599), .ZN(n594) );
  INV_X1 U560 ( .I(n596), .ZN(n599) );
  NOR2_X1 U561 ( .A1(n587), .A2(n588), .ZN(n500) );
  NAND2_X1 U562 ( .A1(activ[4]), .A2(weight[0]), .ZN(n588) );
  NAND2_X1 U563 ( .A1(n600), .A2(n601), .ZN(n587) );
  NAND2_X1 U564 ( .A1(n491), .A2(n602), .ZN(n601) );
  NAND2_X1 U565 ( .A1(n493), .A2(n485), .ZN(n602) );
  INV_X1 U566 ( .I(n488), .ZN(n485) );
  INV_X1 U567 ( .I(n494), .ZN(n491) );
  NAND2_X1 U568 ( .A1(n603), .A2(n604), .ZN(n494) );
  NAND2_X1 U569 ( .A1(n605), .A2(activ[2]), .ZN(n604) );
  NOR2_X1 U570 ( .A1(n606), .A2(n471), .ZN(n605) );
  NOR2_X1 U571 ( .A1(n481), .A2(n475), .ZN(n606) );
  NAND2_X1 U572 ( .A1(n481), .A2(n475), .ZN(n603) );
  NAND2_X1 U573 ( .A1(n607), .A2(n608), .ZN(n475) );
  INV_X1 U574 ( .I(n609), .ZN(n608) );
  NOR2_X1 U575 ( .A1(n610), .A2(n611), .ZN(n609) );
  NAND2_X1 U576 ( .A1(n611), .A2(n610), .ZN(n607) );
  NOR2_X1 U577 ( .A1(n612), .A2(n613), .ZN(n611) );
  NOR2_X1 U578 ( .A1(n610), .A2(n614), .ZN(n481) );
  NAND2_X1 U579 ( .A1(weight[1]), .A2(activ[1]), .ZN(n610) );
  NAND2_X1 U580 ( .A1(n488), .A2(n492), .ZN(n600) );
  INV_X1 U581 ( .I(n493), .ZN(n492) );
  NOR2_X1 U582 ( .A1(n615), .A2(n471), .ZN(n493) );
  INV_X1 U583 ( .I(weight[0]), .ZN(n471) );
  NOR2_X1 U584 ( .A1(n616), .A2(n617), .ZN(n488) );
  INV_X1 U585 ( .I(n618), .ZN(n617) );
  NAND2_X1 U586 ( .A1(n619), .A2(n620), .ZN(n618) );
  NOR2_X1 U587 ( .A1(n620), .A2(n619), .ZN(n616) );
  NOR2_X1 U588 ( .A1(n621), .A2(n622), .ZN(n620) );
  INV_X1 U589 ( .I(n623), .ZN(n622) );
  NAND2_X1 U590 ( .A1(n624), .A2(n625), .ZN(n623) );
  NOR2_X1 U591 ( .A1(n625), .A2(n624), .ZN(n621) );
  NAND2_X1 U592 ( .A1(activ[2]), .A2(weight[1]), .ZN(n625) );
  NOR2_X1 U593 ( .A1(n520), .A2(n526), .ZN(n555) );
  INV_X1 U594 ( .I(n529), .ZN(n526) );
  NOR2_X1 U595 ( .A1(n523), .A2(n529), .ZN(n553) );
  NAND2_X1 U596 ( .A1(activ[7]), .A2(weight[0]), .ZN(n529) );
  INV_X1 U597 ( .I(n520), .ZN(n523) );
  NOR2_X1 U598 ( .A1(n626), .A2(n627), .ZN(n520) );
  NOR2_X1 U599 ( .A1(n628), .A2(n629), .ZN(n627) );
  INV_X1 U600 ( .I(n630), .ZN(n626) );
  NAND2_X1 U601 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U602 ( .A1(n631), .A2(n632), .ZN(n628) );
  NAND2_X1 U603 ( .A1(n633), .A2(n634), .ZN(n632) );
  NOR2_X1 U604 ( .A1(n635), .A2(n534), .ZN(n551) );
  INV_X1 U605 ( .I(n533), .ZN(n534) );
  NOR2_X1 U606 ( .A1(n636), .A2(n637), .ZN(n533) );
  NOR2_X1 U607 ( .A1(n638), .A2(n639), .ZN(n637) );
  INV_X1 U608 ( .I(n640), .ZN(n636) );
  NAND2_X1 U609 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U610 ( .A1(n641), .A2(n642), .ZN(n638) );
  INV_X1 U611 ( .I(n643), .ZN(n639) );
  NOR2_X1 U612 ( .A1(n543), .A2(n544), .ZN(n635) );
  INV_X1 U613 ( .I(n541), .ZN(n543) );
  NAND2_X1 U614 ( .A1(n644), .A2(n645), .ZN(n549) );
  NAND2_X1 U615 ( .A1(n427), .A2(n646), .ZN(n645) );
  INV_X1 U616 ( .I(n429), .ZN(n646) );
  NAND2_X1 U617 ( .A1(n429), .A2(n647), .ZN(n644) );
  INV_X1 U618 ( .I(n427), .ZN(n647) );
  NOR2_X1 U619 ( .A1(n648), .A2(n362), .ZN(n427) );
  INV_X1 U620 ( .I(n369), .ZN(n362) );
  NAND2_X1 U621 ( .A1(n649), .A2(n650), .ZN(n369) );
  NOR2_X1 U622 ( .A1(n650), .A2(n649), .ZN(n648) );
  NOR2_X1 U623 ( .A1(n651), .A2(n652), .ZN(n649) );
  NOR2_X1 U624 ( .A1(n653), .A2(n654), .ZN(n652) );
  INV_X1 U625 ( .I(n422), .ZN(n654) );
  NOR2_X1 U626 ( .A1(n422), .A2(n655), .ZN(n651) );
  INV_X1 U627 ( .I(n653), .ZN(n655) );
  NAND2_X1 U628 ( .A1(n420), .A2(n423), .ZN(n653) );
  NAND2_X1 U629 ( .A1(n656), .A2(n657), .ZN(n423) );
  NAND2_X1 U630 ( .A1(activ[7]), .A2(weight[3]), .ZN(n657) );
  INV_X1 U631 ( .I(n658), .ZN(n656) );
  NAND2_X1 U632 ( .A1(activ[7]), .A2(n658), .ZN(n420) );
  NAND2_X1 U633 ( .A1(n659), .A2(n660), .ZN(n658) );
  NAND2_X1 U634 ( .A1(n661), .A2(n662), .ZN(n660) );
  INV_X1 U635 ( .I(n663), .ZN(n661) );
  NOR2_X1 U636 ( .A1(n664), .A2(n665), .ZN(n422) );
  INV_X1 U637 ( .I(n666), .ZN(n665) );
  NAND2_X1 U638 ( .A1(n417), .A2(n667), .ZN(n666) );
  NOR2_X1 U639 ( .A1(n667), .A2(n417), .ZN(n664) );
  NAND2_X1 U640 ( .A1(n668), .A2(n669), .ZN(n417) );
  NAND2_X1 U641 ( .A1(n670), .A2(n387), .ZN(n669) );
  INV_X1 U642 ( .I(n393), .ZN(n387) );
  INV_X1 U643 ( .I(n671), .ZN(n670) );
  NAND2_X1 U644 ( .A1(n393), .A2(n671), .ZN(n668) );
  NAND2_X1 U645 ( .A1(n672), .A2(n673), .ZN(n671) );
  INV_X1 U646 ( .I(n390), .ZN(n673) );
  NOR2_X1 U647 ( .A1(n388), .A2(n392), .ZN(n390) );
  NAND2_X1 U648 ( .A1(n392), .A2(n674), .ZN(n672) );
  NAND2_X1 U649 ( .A1(weight[5]), .A2(activ[5]), .ZN(n674) );
  NOR2_X1 U650 ( .A1(n675), .A2(n676), .ZN(n392) );
  INV_X1 U651 ( .I(n677), .ZN(n676) );
  NAND2_X1 U652 ( .A1(n678), .A2(n679), .ZN(n677) );
  NAND2_X1 U653 ( .A1(n680), .A2(n681), .ZN(n675) );
  NAND2_X1 U654 ( .A1(n682), .A2(n679), .ZN(n681) );
  NAND2_X1 U655 ( .A1(n683), .A2(n684), .ZN(n393) );
  INV_X1 U656 ( .I(n685), .ZN(n684) );
  NOR2_X1 U657 ( .A1(n401), .A2(n686), .ZN(n685) );
  NAND2_X1 U658 ( .A1(n686), .A2(n401), .ZN(n683) );
  NAND2_X1 U659 ( .A1(n687), .A2(n688), .ZN(n401) );
  NAND2_X1 U660 ( .A1(n689), .A2(n690), .ZN(n688) );
  NAND2_X1 U661 ( .A1(n691), .A2(n692), .ZN(n689) );
  INV_X1 U662 ( .I(n693), .ZN(n687) );
  NOR2_X1 U663 ( .A1(n692), .A2(n691), .ZN(n693) );
  INV_X1 U664 ( .I(n694), .ZN(n691) );
  NAND2_X1 U665 ( .A1(n695), .A2(n696), .ZN(n686) );
  NAND2_X1 U666 ( .A1(n405), .A2(n403), .ZN(n696) );
  NAND2_X1 U667 ( .A1(n404), .A2(n402), .ZN(n695) );
  INV_X1 U668 ( .I(n405), .ZN(n402) );
  NOR2_X1 U669 ( .A1(n408), .A2(n697), .ZN(n405) );
  INV_X1 U670 ( .I(n403), .ZN(n404) );
  NAND2_X1 U671 ( .A1(weight[7]), .A2(activ[3]), .ZN(n403) );
  NOR2_X1 U672 ( .A1(n698), .A2(n699), .ZN(n667) );
  INV_X1 U673 ( .I(n700), .ZN(n699) );
  NAND2_X1 U674 ( .A1(n416), .A2(n418), .ZN(n700) );
  NOR2_X1 U675 ( .A1(n418), .A2(n416), .ZN(n698) );
  NOR2_X1 U676 ( .A1(n701), .A2(n702), .ZN(n416) );
  INV_X1 U677 ( .I(n703), .ZN(n702) );
  NAND2_X1 U678 ( .A1(n704), .A2(n705), .ZN(n703) );
  NAND2_X1 U679 ( .A1(n706), .A2(n707), .ZN(n704) );
  NOR2_X1 U680 ( .A1(n706), .A2(n707), .ZN(n701) );
  NAND2_X1 U681 ( .A1(activ[6]), .A2(weight[4]), .ZN(n418) );
  NAND2_X1 U682 ( .A1(n708), .A2(n709), .ZN(n650) );
  NAND2_X1 U683 ( .A1(n710), .A2(n711), .ZN(n709) );
  NAND2_X1 U684 ( .A1(n712), .A2(n713), .ZN(n710) );
  NAND2_X1 U685 ( .A1(n714), .A2(n715), .ZN(n708) );
  NOR2_X1 U686 ( .A1(n541), .A2(n542), .ZN(n429) );
  INV_X1 U687 ( .I(n544), .ZN(n542) );
  NAND2_X1 U688 ( .A1(n641), .A2(n716), .ZN(n544) );
  NAND2_X1 U689 ( .A1(n643), .A2(n642), .ZN(n716) );
  NAND2_X1 U690 ( .A1(n717), .A2(n718), .ZN(n642) );
  NOR2_X1 U691 ( .A1(n719), .A2(n720), .ZN(n643) );
  INV_X1 U692 ( .I(n721), .ZN(n720) );
  NAND2_X1 U693 ( .A1(n722), .A2(n723), .ZN(n721) );
  NOR2_X1 U694 ( .A1(n723), .A2(n722), .ZN(n719) );
  NOR2_X1 U695 ( .A1(n724), .A2(n725), .ZN(n723) );
  INV_X1 U696 ( .I(n726), .ZN(n725) );
  NAND2_X1 U697 ( .A1(n727), .A2(n728), .ZN(n726) );
  NOR2_X1 U698 ( .A1(n728), .A2(n727), .ZN(n724) );
  INV_X1 U699 ( .I(n729), .ZN(n641) );
  NOR2_X1 U700 ( .A1(n718), .A2(n717), .ZN(n729) );
  NOR2_X1 U701 ( .A1(n730), .A2(n731), .ZN(n717) );
  NOR2_X1 U702 ( .A1(n629), .A2(n634), .ZN(n731) );
  NAND2_X1 U703 ( .A1(n631), .A2(n732), .ZN(n730) );
  INV_X1 U704 ( .I(n733), .ZN(n732) );
  NOR2_X1 U705 ( .A1(n633), .A2(n629), .ZN(n733) );
  NAND2_X1 U706 ( .A1(n734), .A2(n735), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n736), .A2(n737), .ZN(n735) );
  INV_X1 U708 ( .I(n738), .ZN(n734) );
  NOR2_X1 U709 ( .A1(n737), .A2(n736), .ZN(n738) );
  NOR2_X1 U710 ( .A1(n739), .A2(n740), .ZN(n737) );
  NOR2_X1 U711 ( .A1(n741), .A2(n742), .ZN(n740) );
  INV_X1 U712 ( .I(n743), .ZN(n739) );
  NAND2_X1 U713 ( .A1(n742), .A2(n741), .ZN(n743) );
  INV_X1 U714 ( .I(n744), .ZN(n631) );
  NOR2_X1 U715 ( .A1(n634), .A2(n633), .ZN(n744) );
  INV_X1 U716 ( .I(n745), .ZN(n633) );
  NAND2_X1 U717 ( .A1(n746), .A2(n747), .ZN(n745) );
  NAND2_X1 U718 ( .A1(n748), .A2(activ[5]), .ZN(n747) );
  NOR2_X1 U719 ( .A1(n563), .A2(n569), .ZN(n748) );
  NOR2_X1 U720 ( .A1(n566), .A2(n749), .ZN(n746) );
  NOR2_X1 U721 ( .A1(n750), .A2(n563), .ZN(n749) );
  NOR2_X1 U722 ( .A1(n751), .A2(n752), .ZN(n563) );
  NOR2_X1 U723 ( .A1(n753), .A2(n754), .ZN(n752) );
  INV_X1 U724 ( .I(n755), .ZN(n751) );
  NAND2_X1 U725 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U726 ( .A1(n756), .A2(n757), .ZN(n753) );
  NOR2_X1 U727 ( .A1(n388), .A2(n750), .ZN(n566) );
  INV_X1 U728 ( .I(n567), .ZN(n750) );
  NAND2_X1 U729 ( .A1(n758), .A2(n759), .ZN(n567) );
  NAND2_X1 U730 ( .A1(n583), .A2(n760), .ZN(n759) );
  NAND2_X1 U731 ( .A1(n576), .A2(n581), .ZN(n760) );
  NAND2_X1 U732 ( .A1(n761), .A2(n762), .ZN(n583) );
  NAND2_X1 U733 ( .A1(n596), .A2(n763), .ZN(n762) );
  NAND2_X1 U734 ( .A1(n764), .A2(n598), .ZN(n763) );
  INV_X1 U735 ( .I(n592), .ZN(n764) );
  NAND2_X1 U736 ( .A1(n765), .A2(n766), .ZN(n596) );
  NAND2_X1 U737 ( .A1(n767), .A2(activ[2]), .ZN(n766) );
  NOR2_X1 U738 ( .A1(n768), .A2(n569), .ZN(n767) );
  INV_X1 U739 ( .I(weight[1]), .ZN(n569) );
  NOR2_X1 U740 ( .A1(n624), .A2(n619), .ZN(n768) );
  NAND2_X1 U741 ( .A1(n624), .A2(n619), .ZN(n765) );
  NAND2_X1 U742 ( .A1(n769), .A2(n770), .ZN(n619) );
  NAND2_X1 U743 ( .A1(n771), .A2(n772), .ZN(n770) );
  NAND2_X1 U744 ( .A1(n773), .A2(n774), .ZN(n769) );
  INV_X1 U745 ( .I(n772), .ZN(n773) );
  NOR2_X1 U746 ( .A1(n774), .A2(n469), .ZN(n624) );
  NAND2_X1 U747 ( .A1(weight[1]), .A2(activ[0]), .ZN(n469) );
  NAND2_X1 U748 ( .A1(n597), .A2(n592), .ZN(n761) );
  NAND2_X1 U749 ( .A1(n775), .A2(n776), .ZN(n592) );
  NAND2_X1 U750 ( .A1(n777), .A2(n778), .ZN(n776) );
  INV_X1 U751 ( .I(n779), .ZN(n778) );
  NAND2_X1 U752 ( .A1(n779), .A2(n780), .ZN(n775) );
  NAND2_X1 U753 ( .A1(n781), .A2(n782), .ZN(n779) );
  NAND2_X1 U754 ( .A1(n783), .A2(n784), .ZN(n782) );
  NAND2_X1 U755 ( .A1(n785), .A2(n786), .ZN(n781) );
  INV_X1 U756 ( .I(n598), .ZN(n597) );
  NAND2_X1 U757 ( .A1(activ[3]), .A2(weight[1]), .ZN(n598) );
  INV_X1 U758 ( .I(n787), .ZN(n758) );
  NOR2_X1 U759 ( .A1(n581), .A2(n576), .ZN(n787) );
  NOR2_X1 U760 ( .A1(n788), .A2(n789), .ZN(n576) );
  NOR2_X1 U761 ( .A1(n790), .A2(n791), .ZN(n789) );
  INV_X1 U762 ( .I(n792), .ZN(n788) );
  NAND2_X1 U763 ( .A1(n791), .A2(n790), .ZN(n792) );
  NAND2_X1 U764 ( .A1(n793), .A2(n794), .ZN(n790) );
  NAND2_X1 U765 ( .A1(activ[4]), .A2(weight[1]), .ZN(n581) );
  NAND2_X1 U766 ( .A1(activ[6]), .A2(weight[1]), .ZN(n634) );
  NAND2_X1 U767 ( .A1(activ[7]), .A2(weight[1]), .ZN(n718) );
  NOR2_X1 U768 ( .A1(n795), .A2(n796), .ZN(n541) );
  NOR2_X1 U769 ( .A1(n714), .A2(n797), .ZN(n796) );
  INV_X1 U770 ( .I(n712), .ZN(n714) );
  NOR2_X1 U771 ( .A1(n798), .A2(n712), .ZN(n795) );
  NAND2_X1 U772 ( .A1(n799), .A2(n800), .ZN(n712) );
  INV_X1 U773 ( .I(n801), .ZN(n800) );
  NOR2_X1 U774 ( .A1(n802), .A2(n663), .ZN(n801) );
  NAND2_X1 U775 ( .A1(n663), .A2(n802), .ZN(n799) );
  NAND2_X1 U776 ( .A1(n659), .A2(n662), .ZN(n802) );
  NAND2_X1 U777 ( .A1(n803), .A2(n804), .ZN(n662) );
  NAND2_X1 U778 ( .A1(activ[6]), .A2(weight[3]), .ZN(n804) );
  INV_X1 U779 ( .I(n805), .ZN(n803) );
  NAND2_X1 U780 ( .A1(activ[6]), .A2(n805), .ZN(n659) );
  NAND2_X1 U781 ( .A1(n806), .A2(n807), .ZN(n805) );
  NAND2_X1 U782 ( .A1(n808), .A2(n809), .ZN(n807) );
  NAND2_X1 U783 ( .A1(n810), .A2(n811), .ZN(n663) );
  INV_X1 U784 ( .I(n812), .ZN(n811) );
  NOR2_X1 U785 ( .A1(n706), .A2(n813), .ZN(n812) );
  NAND2_X1 U786 ( .A1(n813), .A2(n706), .ZN(n810) );
  NOR2_X1 U787 ( .A1(n814), .A2(n815), .ZN(n706) );
  INV_X1 U788 ( .I(n816), .ZN(n815) );
  NAND2_X1 U789 ( .A1(n817), .A2(n679), .ZN(n816) );
  NOR2_X1 U790 ( .A1(n679), .A2(n817), .ZN(n814) );
  NOR2_X1 U791 ( .A1(n818), .A2(n819), .ZN(n817) );
  INV_X1 U792 ( .I(n680), .ZN(n819) );
  NAND2_X1 U793 ( .A1(activ[4]), .A2(n682), .ZN(n680) );
  NOR2_X1 U794 ( .A1(n682), .A2(n678), .ZN(n818) );
  NOR2_X1 U795 ( .A1(n697), .A2(n389), .ZN(n678) );
  INV_X1 U796 ( .I(activ[4]), .ZN(n697) );
  NAND2_X1 U797 ( .A1(n820), .A2(n821), .ZN(n682) );
  NAND2_X1 U798 ( .A1(n822), .A2(n823), .ZN(n821) );
  NAND2_X1 U799 ( .A1(n824), .A2(n825), .ZN(n823) );
  INV_X1 U800 ( .I(n826), .ZN(n820) );
  NOR2_X1 U801 ( .A1(n825), .A2(n824), .ZN(n826) );
  INV_X1 U802 ( .I(n827), .ZN(n825) );
  NOR2_X1 U803 ( .A1(n828), .A2(n829), .ZN(n679) );
  NOR2_X1 U804 ( .A1(n830), .A2(n692), .ZN(n829) );
  INV_X1 U805 ( .I(n831), .ZN(n828) );
  NAND2_X1 U806 ( .A1(n830), .A2(n692), .ZN(n831) );
  NAND2_X1 U807 ( .A1(weight[6]), .A2(activ[3]), .ZN(n692) );
  NAND2_X1 U808 ( .A1(n832), .A2(n833), .ZN(n830) );
  INV_X1 U809 ( .I(n834), .ZN(n833) );
  NOR2_X1 U810 ( .A1(n690), .A2(n694), .ZN(n834) );
  NAND2_X1 U811 ( .A1(n694), .A2(n690), .ZN(n832) );
  NAND2_X1 U812 ( .A1(n835), .A2(n836), .ZN(n690) );
  NAND2_X1 U813 ( .A1(n694), .A2(n837), .ZN(n835) );
  NOR2_X1 U814 ( .A1(n838), .A2(n839), .ZN(n694) );
  NAND2_X1 U815 ( .A1(n840), .A2(n841), .ZN(n813) );
  INV_X1 U816 ( .I(n842), .ZN(n841) );
  NOR2_X1 U817 ( .A1(n705), .A2(n707), .ZN(n842) );
  NAND2_X1 U818 ( .A1(n707), .A2(n705), .ZN(n840) );
  NAND2_X1 U819 ( .A1(n843), .A2(n844), .ZN(n705) );
  NAND2_X1 U820 ( .A1(n845), .A2(n846), .ZN(n844) );
  NAND2_X1 U821 ( .A1(n847), .A2(n848), .ZN(n845) );
  NAND2_X1 U822 ( .A1(n849), .A2(n850), .ZN(n843) );
  NOR2_X1 U823 ( .A1(n388), .A2(n851), .ZN(n707) );
  INV_X1 U824 ( .I(n797), .ZN(n798) );
  NAND2_X1 U825 ( .A1(n852), .A2(n853), .ZN(n797) );
  INV_X1 U826 ( .I(n854), .ZN(n853) );
  NOR2_X1 U827 ( .A1(n711), .A2(n715), .ZN(n854) );
  NAND2_X1 U828 ( .A1(n715), .A2(n711), .ZN(n852) );
  NAND2_X1 U829 ( .A1(n855), .A2(n856), .ZN(n711) );
  NAND2_X1 U830 ( .A1(n727), .A2(n857), .ZN(n856) );
  NAND2_X1 U831 ( .A1(n722), .A2(n728), .ZN(n857) );
  NOR2_X1 U832 ( .A1(n858), .A2(n859), .ZN(n727) );
  NOR2_X1 U833 ( .A1(n741), .A2(n860), .ZN(n859) );
  INV_X1 U834 ( .I(n861), .ZN(n860) );
  NAND2_X1 U835 ( .A1(n742), .A2(n736), .ZN(n861) );
  NAND2_X1 U836 ( .A1(n756), .A2(n862), .ZN(n741) );
  NAND2_X1 U837 ( .A1(n754), .A2(n757), .ZN(n862) );
  NAND2_X1 U838 ( .A1(n863), .A2(n864), .ZN(n757) );
  NAND2_X1 U839 ( .A1(activ[4]), .A2(weight[2]), .ZN(n864) );
  INV_X1 U840 ( .I(n865), .ZN(n863) );
  NAND2_X1 U841 ( .A1(n866), .A2(n867), .ZN(n754) );
  INV_X1 U842 ( .I(n868), .ZN(n867) );
  NOR2_X1 U843 ( .A1(n869), .A2(n870), .ZN(n868) );
  NAND2_X1 U844 ( .A1(n870), .A2(n869), .ZN(n866) );
  NAND2_X1 U845 ( .A1(n871), .A2(n872), .ZN(n869) );
  NAND2_X1 U846 ( .A1(activ[4]), .A2(n865), .ZN(n756) );
  NAND2_X1 U847 ( .A1(n793), .A2(n873), .ZN(n865) );
  NAND2_X1 U848 ( .A1(n791), .A2(n794), .ZN(n873) );
  NAND2_X1 U849 ( .A1(n874), .A2(n875), .ZN(n794) );
  NAND2_X1 U850 ( .A1(activ[3]), .A2(weight[2]), .ZN(n875) );
  INV_X1 U851 ( .I(n876), .ZN(n874) );
  NAND2_X1 U852 ( .A1(n877), .A2(n878), .ZN(n791) );
  NAND2_X1 U853 ( .A1(n879), .A2(n880), .ZN(n878) );
  INV_X1 U854 ( .I(n881), .ZN(n877) );
  NOR2_X1 U855 ( .A1(n880), .A2(n879), .ZN(n881) );
  NOR2_X1 U856 ( .A1(n882), .A2(n883), .ZN(n880) );
  INV_X1 U857 ( .I(n884), .ZN(n883) );
  NAND2_X1 U858 ( .A1(n885), .A2(n886), .ZN(n884) );
  NOR2_X1 U859 ( .A1(n886), .A2(n885), .ZN(n882) );
  NAND2_X1 U860 ( .A1(weight[3]), .A2(activ[2]), .ZN(n886) );
  NAND2_X1 U861 ( .A1(activ[3]), .A2(n876), .ZN(n793) );
  NAND2_X1 U862 ( .A1(n887), .A2(n888), .ZN(n876) );
  NAND2_X1 U863 ( .A1(n777), .A2(n889), .ZN(n888) );
  NAND2_X1 U864 ( .A1(n786), .A2(n784), .ZN(n889) );
  INV_X1 U865 ( .I(n785), .ZN(n784) );
  INV_X1 U866 ( .I(n783), .ZN(n786) );
  INV_X1 U867 ( .I(n780), .ZN(n777) );
  NOR2_X1 U868 ( .A1(n890), .A2(n891), .ZN(n780) );
  NOR2_X1 U869 ( .A1(n892), .A2(n893), .ZN(n891) );
  INV_X1 U870 ( .I(n894), .ZN(n890) );
  NAND2_X1 U871 ( .A1(n893), .A2(n892), .ZN(n894) );
  NAND2_X1 U872 ( .A1(weight[3]), .A2(activ[1]), .ZN(n892) );
  INV_X1 U873 ( .I(n895), .ZN(n893) );
  NAND2_X1 U874 ( .A1(n785), .A2(n783), .ZN(n887) );
  NOR2_X1 U875 ( .A1(n839), .A2(n612), .ZN(n783) );
  NOR2_X1 U876 ( .A1(n772), .A2(n774), .ZN(n785) );
  INV_X1 U877 ( .I(n771), .ZN(n774) );
  NOR2_X1 U878 ( .A1(n612), .A2(n470), .ZN(n771) );
  NOR2_X1 U879 ( .A1(n736), .A2(n742), .ZN(n858) );
  NOR2_X1 U880 ( .A1(n388), .A2(n612), .ZN(n742) );
  INV_X1 U881 ( .I(weight[2]), .ZN(n612) );
  INV_X1 U882 ( .I(activ[5]), .ZN(n388) );
  NAND2_X1 U883 ( .A1(n896), .A2(n897), .ZN(n736) );
  INV_X1 U884 ( .I(n898), .ZN(n897) );
  NOR2_X1 U885 ( .A1(n899), .A2(n900), .ZN(n898) );
  NAND2_X1 U886 ( .A1(n900), .A2(n899), .ZN(n896) );
  NAND2_X1 U887 ( .A1(n901), .A2(n902), .ZN(n899) );
  INV_X1 U888 ( .I(n903), .ZN(n855) );
  NOR2_X1 U889 ( .A1(n722), .A2(n728), .ZN(n903) );
  NAND2_X1 U890 ( .A1(activ[6]), .A2(weight[2]), .ZN(n728) );
  NAND2_X1 U891 ( .A1(n904), .A2(n905), .ZN(n722) );
  NAND2_X1 U892 ( .A1(n906), .A2(n808), .ZN(n905) );
  INV_X1 U893 ( .I(n907), .ZN(n906) );
  NAND2_X1 U894 ( .A1(n908), .A2(n907), .ZN(n904) );
  NAND2_X1 U895 ( .A1(n806), .A2(n809), .ZN(n907) );
  NAND2_X1 U896 ( .A1(n909), .A2(n910), .ZN(n809) );
  NAND2_X1 U897 ( .A1(activ[5]), .A2(weight[3]), .ZN(n910) );
  INV_X1 U898 ( .I(n911), .ZN(n909) );
  NAND2_X1 U899 ( .A1(activ[5]), .A2(n911), .ZN(n806) );
  NAND2_X1 U900 ( .A1(n901), .A2(n912), .ZN(n911) );
  NAND2_X1 U901 ( .A1(n900), .A2(n902), .ZN(n912) );
  NAND2_X1 U902 ( .A1(n913), .A2(n914), .ZN(n902) );
  NAND2_X1 U903 ( .A1(activ[4]), .A2(weight[3]), .ZN(n914) );
  INV_X1 U904 ( .I(n915), .ZN(n913) );
  NAND2_X1 U905 ( .A1(n916), .A2(n917), .ZN(n900) );
  NAND2_X1 U906 ( .A1(n918), .A2(n919), .ZN(n917) );
  INV_X1 U907 ( .I(n920), .ZN(n916) );
  NOR2_X1 U908 ( .A1(n919), .A2(n918), .ZN(n920) );
  NOR2_X1 U909 ( .A1(n921), .A2(n922), .ZN(n919) );
  NOR2_X1 U910 ( .A1(n923), .A2(n924), .ZN(n922) );
  INV_X1 U911 ( .I(n925), .ZN(n921) );
  NAND2_X1 U912 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U913 ( .A1(activ[4]), .A2(n915), .ZN(n901) );
  NAND2_X1 U914 ( .A1(n871), .A2(n926), .ZN(n915) );
  NAND2_X1 U915 ( .A1(n870), .A2(n872), .ZN(n926) );
  NAND2_X1 U916 ( .A1(n927), .A2(n928), .ZN(n872) );
  NAND2_X1 U917 ( .A1(activ[3]), .A2(weight[3]), .ZN(n928) );
  INV_X1 U918 ( .I(n929), .ZN(n927) );
  NAND2_X1 U919 ( .A1(n930), .A2(n931), .ZN(n870) );
  INV_X1 U920 ( .I(n932), .ZN(n931) );
  NOR2_X1 U921 ( .A1(n933), .A2(n934), .ZN(n932) );
  NAND2_X1 U922 ( .A1(n934), .A2(n933), .ZN(n930) );
  NAND2_X1 U923 ( .A1(n935), .A2(n936), .ZN(n934) );
  NAND2_X1 U924 ( .A1(n937), .A2(n938), .ZN(n936) );
  INV_X1 U925 ( .I(n939), .ZN(n935) );
  NOR2_X1 U926 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U927 ( .A1(activ[3]), .A2(n929), .ZN(n871) );
  NAND2_X1 U928 ( .A1(n940), .A2(n941), .ZN(n929) );
  NAND2_X1 U929 ( .A1(n942), .A2(weight[3]), .ZN(n941) );
  NOR2_X1 U930 ( .A1(n943), .A2(n839), .ZN(n942) );
  NOR2_X1 U931 ( .A1(n885), .A2(n879), .ZN(n943) );
  NAND2_X1 U932 ( .A1(n885), .A2(n879), .ZN(n940) );
  NAND2_X1 U933 ( .A1(n944), .A2(n945), .ZN(n879) );
  INV_X1 U934 ( .I(n946), .ZN(n945) );
  NOR2_X1 U935 ( .A1(n947), .A2(n948), .ZN(n946) );
  NAND2_X1 U936 ( .A1(n948), .A2(n947), .ZN(n944) );
  NOR2_X1 U937 ( .A1(n947), .A2(n772), .ZN(n885) );
  NAND2_X1 U938 ( .A1(weight[3]), .A2(activ[0]), .ZN(n772) );
  NAND2_X1 U939 ( .A1(weight[4]), .A2(activ[1]), .ZN(n947) );
  INV_X1 U940 ( .I(n808), .ZN(n908) );
  NOR2_X1 U941 ( .A1(n949), .A2(n950), .ZN(n808) );
  NOR2_X1 U942 ( .A1(n847), .A2(n951), .ZN(n950) );
  INV_X1 U943 ( .I(n952), .ZN(n949) );
  NAND2_X1 U944 ( .A1(n951), .A2(n847), .ZN(n952) );
  INV_X1 U945 ( .I(n849), .ZN(n847) );
  NAND2_X1 U946 ( .A1(n953), .A2(n954), .ZN(n849) );
  INV_X1 U947 ( .I(n955), .ZN(n954) );
  NOR2_X1 U948 ( .A1(n824), .A2(n956), .ZN(n955) );
  NAND2_X1 U949 ( .A1(n956), .A2(n824), .ZN(n953) );
  NOR2_X1 U950 ( .A1(n957), .A2(n958), .ZN(n824) );
  INV_X1 U951 ( .I(n959), .ZN(n958) );
  NAND2_X1 U952 ( .A1(n960), .A2(n961), .ZN(n959) );
  NOR2_X1 U953 ( .A1(n961), .A2(n960), .ZN(n957) );
  NOR2_X1 U954 ( .A1(n408), .A2(n839), .ZN(n960) );
  NAND2_X1 U955 ( .A1(n962), .A2(n836), .ZN(n961) );
  NAND2_X1 U956 ( .A1(n962), .A2(n963), .ZN(n836) );
  NOR2_X1 U957 ( .A1(n838), .A2(n470), .ZN(n962) );
  INV_X1 U958 ( .I(weight[7]), .ZN(n838) );
  NAND2_X1 U959 ( .A1(n964), .A2(n965), .ZN(n956) );
  INV_X1 U960 ( .I(n966), .ZN(n965) );
  NOR2_X1 U961 ( .A1(n822), .A2(n827), .ZN(n966) );
  NAND2_X1 U962 ( .A1(n827), .A2(n822), .ZN(n964) );
  NAND2_X1 U963 ( .A1(n967), .A2(n968), .ZN(n822) );
  NAND2_X1 U964 ( .A1(n969), .A2(weight[5]), .ZN(n968) );
  NOR2_X1 U965 ( .A1(n970), .A2(n839), .ZN(n969) );
  INV_X1 U966 ( .I(activ[2]), .ZN(n839) );
  NOR2_X1 U967 ( .A1(n971), .A2(n972), .ZN(n970) );
  NAND2_X1 U968 ( .A1(n971), .A2(n972), .ZN(n967) );
  NOR2_X1 U969 ( .A1(n389), .A2(n615), .ZN(n827) );
  NAND2_X1 U970 ( .A1(n973), .A2(n974), .ZN(n951) );
  NAND2_X1 U971 ( .A1(n975), .A2(n850), .ZN(n974) );
  NAND2_X1 U972 ( .A1(n848), .A2(n846), .ZN(n973) );
  INV_X1 U973 ( .I(n975), .ZN(n846) );
  NOR2_X1 U974 ( .A1(n976), .A2(n977), .ZN(n975) );
  INV_X1 U975 ( .I(n978), .ZN(n977) );
  NAND2_X1 U976 ( .A1(n979), .A2(n923), .ZN(n978) );
  NAND2_X1 U977 ( .A1(n980), .A2(n981), .ZN(n923) );
  INV_X1 U978 ( .I(n982), .ZN(n981) );
  NOR2_X1 U979 ( .A1(n983), .A2(n937), .ZN(n982) );
  NOR2_X1 U980 ( .A1(n984), .A2(n895), .ZN(n937) );
  NAND2_X1 U981 ( .A1(weight[4]), .A2(activ[0]), .ZN(n895) );
  NOR2_X1 U982 ( .A1(n938), .A2(n933), .ZN(n983) );
  NAND2_X1 U983 ( .A1(n933), .A2(n938), .ZN(n980) );
  NAND2_X1 U984 ( .A1(weight[4]), .A2(activ[2]), .ZN(n938) );
  NOR2_X1 U985 ( .A1(n985), .A2(n986), .ZN(n933) );
  NOR2_X1 U986 ( .A1(n984), .A2(n963), .ZN(n986) );
  INV_X1 U987 ( .I(n987), .ZN(n985) );
  NAND2_X1 U988 ( .A1(n963), .A2(n984), .ZN(n987) );
  NAND2_X1 U989 ( .A1(weight[5]), .A2(activ[1]), .ZN(n984) );
  NOR2_X1 U990 ( .A1(n408), .A2(n613), .ZN(n963) );
  NAND2_X1 U991 ( .A1(n924), .A2(n918), .ZN(n979) );
  NOR2_X1 U992 ( .A1(n918), .A2(n924), .ZN(n976) );
  NOR2_X1 U993 ( .A1(n851), .A2(n615), .ZN(n924) );
  INV_X1 U994 ( .I(activ[3]), .ZN(n615) );
  INV_X1 U995 ( .I(weight[4]), .ZN(n851) );
  NAND2_X1 U996 ( .A1(n988), .A2(n989), .ZN(n918) );
  NAND2_X1 U997 ( .A1(n972), .A2(n990), .ZN(n989) );
  INV_X1 U998 ( .I(n991), .ZN(n988) );
  NOR2_X1 U999 ( .A1(n990), .A2(n972), .ZN(n991) );
  NAND2_X1 U1000 ( .A1(n992), .A2(n993), .ZN(n972) );
  NAND2_X1 U1001 ( .A1(n837), .A2(n994), .ZN(n993) );
  INV_X1 U1002 ( .I(n995), .ZN(n992) );
  NOR2_X1 U1003 ( .A1(n994), .A2(n837), .ZN(n995) );
  NAND2_X1 U1004 ( .A1(weight[7]), .A2(activ[0]), .ZN(n994) );
  NOR2_X1 U1005 ( .A1(n996), .A2(n997), .ZN(n990) );
  NOR2_X1 U1006 ( .A1(n998), .A2(n999), .ZN(n997) );
  INV_X1 U1007 ( .I(n1000), .ZN(n999) );
  NOR2_X1 U1008 ( .A1(n1000), .A2(n971), .ZN(n996) );
  INV_X1 U1009 ( .I(n998), .ZN(n971) );
  NAND2_X1 U1010 ( .A1(n837), .A2(n948), .ZN(n998) );
  NOR2_X1 U1011 ( .A1(n389), .A2(n613), .ZN(n948) );
  INV_X1 U1012 ( .I(activ[0]), .ZN(n613) );
  INV_X1 U1013 ( .I(weight[5]), .ZN(n389) );
  NOR2_X1 U1014 ( .A1(n408), .A2(n470), .ZN(n837) );
  INV_X1 U1015 ( .I(activ[1]), .ZN(n470) );
  INV_X1 U1016 ( .I(weight[6]), .ZN(n408) );
  NAND2_X1 U1017 ( .A1(weight[5]), .A2(activ[2]), .ZN(n1000) );
  INV_X1 U1018 ( .I(n850), .ZN(n848) );
  NAND2_X1 U1019 ( .A1(weight[4]), .A2(activ[4]), .ZN(n850) );
  INV_X1 U1020 ( .I(n713), .ZN(n715) );
  NAND2_X1 U1021 ( .A1(activ[7]), .A2(weight[2]), .ZN(n713) );
  NAND2_X1 U1022 ( .A1(n1001), .A2(n1002), .ZN(out[0]) );
  NAND2_X1 U1023 ( .A1(prev_mac_o[0]), .A2(n614), .ZN(n1002) );
  NAND2_X1 U1024 ( .A1(n472), .A2(n1003), .ZN(n1001) );
  INV_X1 U1025 ( .I(prev_mac_o[0]), .ZN(n1003) );
  INV_X1 U1026 ( .I(n614), .ZN(n472) );
  NAND2_X1 U1027 ( .A1(weight[0]), .A2(activ[0]), .ZN(n614) );
endmodule

